module klingon_dataf(
  input [3:0] I,
  output [6:0] O
);

  wire [3:0] i;
  assign i = I[3:0];

  assign O = (i == 0) ? 7'b1111110 :
             (i == 1) ? 7'b1000000 :
             (i == 2) ? 7'b1000001 :
             (i == 3) ? 7'b1001001 :
             (i == 4) ? 7'b0100011 :
             (i == 5) ? 7'b0011101 :
             (i == 6) ? 7'b0100101 :
             (i == 7) ? 7'b0000111 :
             (i == 8) ? 7'b0100111 :
             (i == 9) ? 7'b0101111 :
             7'b0000000;

endmodule
